* VREG *
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include ../schem/voltage-reg.spice

.param pvdd=5.0V
.param pvss=0.0V
.param pvb1=5.0V
.param pvb2=1.7V

Vdd VDD GND SIN('pvdd' 10mV 100KHz)
Vss VSS GND DC 'pvss'
Vb1 VB1 GND DC 'pvb1'
Vb2 VB2 GND DC 'pvb2'
*Vnoise VDD V SIN(0 1m 10KHz)

*.noise v(OUT) Vdd dec 10 1kHz 100MEG

Xreg OUT VB2 VB1 voltage-reg

.control
tran 0.1m 20m 0m
*noise v(OUT) Vdd dec 10 1kHz 100MEG
plot V(OUT)
plot V(VDD)

.endc


.end
