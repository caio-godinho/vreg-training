* VREG *
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include ../schem/voltage-reg.spice

.param pvdd=5.0V
.param pvss=0.0V
.param pvb1=5.0V
.param pvb2=1.7V
*.param pcap=0.0pF
.param pres=0.0KOhm

Vdd VDD GND SIN('pvdd' 10mV 100KHz)
Vss VSS GND DC 'pvss'
Vb1 VB1 GND DC 'pvb1'
Vb2 VB2 GND DC 'pvb2'

Xreg OUT VB2 VB1 voltage-reg

*Cout OUT GND 'pcap'
Rout OUT GND 'pres'

**.include control-commands/capacitiveLoad-var.spice
.include control-commands/resistiveLoad-var.spice


.end
