** sch_path: /home/caio-godinho/repos/vreg-training/schem/voltage-reg.sch
.subckt voltage-reg OUT VB2 VB1
*.PININFO OUT:O VB2:I VB1:I
XM1 VDD VB1 OUT GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=1
XM2 VSS VB2 OUT VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W='7*2.8125' nf=1 m=1
.ends
.GLOBAL VDD
.GLOBAL VSS
.GLOBAL GND
.end
